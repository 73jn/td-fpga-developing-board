.SUBCKT MCP651 1 2 3 4 5
*              | | | | |
*              | | | | Output
*              | | | Negative Supply
*              | | Positive Supply
*              | Inverting Input
*              Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP651, MCP652, MCP655
*
* Revision History:
*      REV A: 26-Oct-09, Created model
*       
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*      If you have a problem with your circuit, make sure to check the input
*      terminal voltages against the common mode input range.
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Some Variation in specs vs. Power Supply Voltage
*      Vos distribution, Ib distribution for Monte Carlo
*      Distortion (detailed non-linear behavior)
*      Some Temperature analysis
*      Process variation
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 -500M
R10 10 11 100k
R11 10 12 100k
G10 10 11 10 11 10M
G11 10 12 10 12 10M
C12  1  0 9.00P
E12 71 14 POLY(4) 205 0 222 0 26 0 27 0 200U 54 1.27 1 1
G12 1 0 62 0 1m
G13 1 2 63 0 1u
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 1m
C14  2  0 9.00P
I15 15 4 1
V16 16 4 -.3
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 1.3
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 12E12
R72  2  0 12E12
R73  1  2 20E12
*
* Noise, PSRR, and CMRR
I20 21 20 423u
D20 20  0 DN1
D21  0 21 DN1
E21 201 0 POLY(2) 20 0 21 0 0 1 1
R201 201 204 .5
C201 204 202 100u
R202 202 0   30m
R203 203 0   18m
C203 202 203 2.5m
R204 204 205 4
C204 204 205 50u
C205 205 206 50u
R205 206 0  .5
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
E22 221 0 POLY(2) 22 0 23 0 0 1 1
R221 221 222 1
C221 222 0 93n
G26  0 26 POLY(2) 3 0 4 0   0.00 -56.2U -56.2U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -.37M 79U 79U
R27 27 0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 4.36
I31 0 31 DC 13.5
R31 31  0 1 TC=1.8M,-5U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 3.94
I32 32 0 DC 21.1
R32 32  0 1 TC=1.35M,-5U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
C33 33 0 1.6p
G34  0 34 33 0 1
R34  34 0 1K
C34  34 0 0.72U
G38  0 38 34 0 100m
R38  39 0 10
L38  38 39 7N
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(0.64,1n))(0.65,2))
G36 33 0 TABLE {V(35,4)} ((-1.46,-1)((-1.45,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57 0 25
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0 0 12.5M 2.3M 33.3M
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
CD55 55 57 2p
CD56 57 56 2p
E55 55  0 POLY(3) 3 0 51 0 3 4 -3.1M 1 -4.6M 4M 0 0 -0m 0 -0.5m
E56 56  0 POLY(3) 4 0 52 0 3 4 1.7M 1 -6.7M 0M 0 0 0m 0 -0.28m
**                       0 3 4 -lowend-same 1 mainR divergLow 0 0 hiDiff 0 sl_fn(isq)
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -1 1M
G54  0  4 POLY(1) 52 0  -1 -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-173U,-199N
G97 0 98 TABLE { V(96,5) } ((-11,-96M)(-1M,-95M)(0,0)(1M,95M)(11,96M))
E97 99 0 VALUE { V(98)*((V(3)-V(4))*-6.72M + 1.01)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=2.78M,2.41U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(1.2,1u)(1.3,54.0U)(1.5,500U)(1.8,4.3M)
+ (2.5,5.00M)(3.5,5.4M)(6.5,6.1M))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=2.5
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 REXP  2.5M
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1uA
R63 0 63 5.00 TC=-3M,0.8M
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L & W values
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=146E-18 AF=1
.MODEL REXP  RES TCE= 6.7
.ENDS MCP651
