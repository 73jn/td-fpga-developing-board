.SUBCKT MCP6051 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP6051, MCP6052, MCP6054
*
* Revision History:
*      REV A: 19-Aug-09, Created model
*
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Some Variation in specs vs. Power Supply Voltage
*      Vos distribution, Ib distribution for Monte Carlo
*      Distortion (detailed non-linear behavior)
*      Some Temperature analysis
*      Process variation
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 -500M
R10 10 11 2.18MEG
R11 10 12 2.18MEG
G10 10 11 10 11 40U
G11 10 12 10 12 40U
C11 11 12 364E-15
C12  1  0 6P
E12 71 14 POLY(6) 20 0 21 0 22 0 23 0 26 0 27 0 100U 13 13 4.7 4.7 1 1
G12 1 0 62 0 1m
G13 1 2 63 0 1u
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 1m
C14  2  0 6P
C13  1  2 3P
I15 15 4 5.00U
V16 16 4 -300M
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 -300M
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 13.3E12
R72  2  0 13.3E12
R73  1  2 13.3E12
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G26  0 26 POLY(2) 3 0 4 0   0.00 -63.0U -8.91U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -2120N 100N 100N
R27 27 0 0.1m
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 6.5
I31 0 31 DC 43
R31 31  0 1 TC=3.0M,-1U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 4
I32 32 0 DC 80
R32 32  0 1 TC=2.4M,-6U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 562M
R34  34 0 1K
C34  34 0 235U
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 88.4P
G38  0 38 37 0 1m
R38  38 0 1K
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(270,1n))(297,1))
G36 33 0 TABLE {V(35,4)} ((-297,-1)((-270,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 1.8K
C58  5  0 2.00P
G57  0 57 POLY(4) 3 0 4 0 35 0 27 0 0 0.3M 0.25M 555U .5
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
E55 55  0 POLY(3) 3 0 51 0 3 4 -7M  1 -70.7M -2.2M 0 0 0.56m  0 6.4m
E56 56  0 POLY(3) 4 0 52 0 3 4 6M 1 -60.0M 2M 0 0 0.513m 0 5m
**                   0 3 4 lowend-same 1 mainR divergLow 0 0 hiDiff
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -5.00U 1M
G54  0  4 POLY(1) 52 0  -5.00U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-5.4M,20.3U
G97 0 98 TABLE { V(96,5) } ((-12.0,-7.5m)(-1.00M,-7.42m)(0,0)(1.00M,7.42m)(12.0,7.5m))
E97 99 0 VALUE { V(98)*((V(3)-V(4))*650M + -300M)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=3.05M,-10.0U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(600M,320N)(700M,1.2U)(1.3,26.0U)
+ (1.4,27.0U)(5.2,32.0U)(7.00,34.0U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=1.75,8M
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 REXP 0.9M
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1uA
R63 0 63 950M TC=6M,0.52M
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L & W values
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=146E-18 AF=1
.MODEL REXP  RES TCE= 7.2
.ENDS MCP6051
