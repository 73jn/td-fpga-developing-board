.SUBCKT MCP6071 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP6071, MCP6072, MCP6074
*
* Revision History:
*      REV A: 03-Aug-09, Created model
*      
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Some Variation in specs vs. Power Supply Voltage
*      Vos distribution, Ib distribution for Monte Carlo
*      Distortion (detailed non-linear behavior)
*      Common Mode Input Range does not vary with Vdd in model, use Fig 2-13 for critical apps
*      Some Temperature analysis
*      Process variation
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 -500M
R10 10 11 500k
R11 10 12 500k
G10 10 11 10 11 0.215M
G11 10 12 10 12 0.215M
C11 11 12 165P
C12  1  0 6P
C13  1  2 3P
E12 71 14 POLY(4) 20 0 21 0 26 0 27 0 160U 14.7 14.7 1 1
G12 1 0 62 0 1m
G13 1 2 63 0 1u
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 1m
C14  2  0 6P
I15 15 4 100U
V16 16 4 -300M
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 -300M
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 20.0E12
R72  2  0 20.0E12
R73  1  2 20.0E12
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
G26  0 26 POLY(2) 3 0 4 0   0.00 -70U -7.5U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -138U 9U 9U
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 5
I31 0 31 DC 40
R31 31  0 1 TC=2.76M,-14.3U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 0.45
I32 32 0 DC 85
R32 32  0 1 TC=2.75M,-14.3U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 562M
R34  34 0 1K
C34  34 0 70U
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 40P
G38  0 38 37 0 1m
R38  39 0 1K
L38  38 39 1.6M
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(61,1n))(62,1))
G36 33 0 TABLE {V(35,4)} ((-61,-1)((-60,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 500
*R57 57  0 250
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0   0 2M 0.82M 2M
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G55 0 551 POLY(2) 3 0 51 0 -.99M 1 -32M
G56 0 561 POLY(2) 4 0 52 0 1.14M 1 -29M
R55 551 0 1 TC=-12U
R56 561 0 1 TC=-15U, -30N
E55 55 0 551 0 1
E56 56 0 561 0 1
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -100U 1M
G54  0  4 POLY(1) 52 0  -100U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-4.8M,22U
G97 0 98 TABLE {V(96,5)} ((-11,-10.1M)(-1M,-10M)(0,0)(1M,10M)(11,10.1M))
E97 99 0 VALUE {V(98)*((V(3)-V(4))*470M + -40M)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=3M
G61 3 4 61 0 1
G60 0 61 TABLE {V(3,4)} 
+ ((0,0)(900M,10N)(1,15U)(1.4,96U)(1.5,99U)(7,118U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=-0.5, -60m
E75 1 71 70 0 1
*
* Temp Sensistive IBias
I62 0 62 DC 1UA
R62 0 621 REXP  300U
R621 621 62 RLIN 0.6M
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1uA
R63 0 63 0.97 TC=2.5M,0.62M
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L & W values
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=146E-18 AF=1
.MODEL REXP  RES TCE= 8.4
.MODEL RLIN	 RES TC1= .15 TC2= 2M  
.ENDS MCP6071
