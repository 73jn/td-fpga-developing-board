.SUBCKT MCP6285 1 2 3 4 5 6 7
*               | | | | | | |
*               | | | | | | Output Amp 2
*               | | | | | Inverting Input Amp 2 
*               | | | | Output Amp 1/Non-inverting Input Amp 2
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input amp 1
*               Non-inverting Input amp 1
X1 1 2 3 4 5 MCP6281
X2 5 6 3 4 7 MCP6281
.ENDS
*
.SUBCKT MCP6281 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP6281,MCP6282,MCP6283,MCP6284,MCP6285
*
* Revision History:
*      REV A: 23-Aug-06, HNV (created model)  
*	                     (MC_RP, 23-Aug-06, Level 1.16)
*       
* Recommendations:
*      Use PSPICE (other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Chip select (MCP6283, MCP6285)
*      Some Variation in specs vs. Power Supply Voltage
*      Monte Carlo (Vos, Ib), Process variation
*      Distortion (detailed non-linear behavior)
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 -500M
R10 10 11 1MEG
R11 10 12 1MEG
G10 10 11 10 11 150u
G11 10 12 10 12 150u
C11 11 12 0.75P
C12  1  0 6.00P
E12 71 14 POLY(4) 20 0 21 0 26 0 27 0   3.00M 7 7 1 1
G12 1 0 62 0 1m
M12 11 14 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G13 1 2 62 0 .42m
M14 12 2 15 15 NMI L=2.00U W=42.0U; *Added L & W values
G14 2 0 62 0 1m
C14  2  0 6.00P
I15 15 4 50.0U
V16 16 4 -300M
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 -300M
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 20.0E12
R72  2  0 20.0E12
R73  1  2 20.0E12
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
G26  0 26 POLY(2) 3 0 4 0   0.00 10U 13U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -82.2U 4U 4U
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 -4.77
I31 0 31 DC 97.1
R31 31  0 1 TC=3.44M,1.20U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,.1)(2m,2))
G32 32 0 3 4 -5.94
I32 32 0 DC 121
R32 32  0 1 TC=2.45M,-3.91U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 316M
R34  34 0 1K
C34  34 0 9.4U
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 1.3P
G38  0 38 37 0 1m
R38  39 0 1K
L38  38 39 32U
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(60,1n))(61,1))
G36 33 0 TABLE {V(35,4)} ((-61,-1)((-60,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 500
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0   0 16M 16M 2.00M
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
E55 55  0 POLY(2) 3 0 51 0 -1.2M 1 -20M
E56 56  0 POLY(2) 4 0 52 0 1.4M 1 -18M
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -50.0U 1M
G54  0  4 POLY(1) 52 0  -50.0U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=2.16M,-4.76U
G97 0 98 TABLE { V(96,5) } ((-11.0,-24.0M)(-1.00M,-23.7M)(0,0)(1.00M,23.7M)(11.0,24.0M))
E97 99 0 VALUE { V(98)*((V(3)-V(4))*-66.6M + 1.2)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=2.38M,-3.46U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(800M,4.00U)(950M,20.0U)(1.7,380U)
+ (1.8,390U)(2.00,400U)(5.5,436U))
*
* Temperature Sensistive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=1.7
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 REXP  237.67473U
*
* Models
.MODEL NMI NMOS(KP=20.0U LEVEL=1 ); *Removed L & W values
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=1F AF=1
.MODEL REXP RES TCE= 9.26823
.ENDS MCP6281
