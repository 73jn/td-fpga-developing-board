--
-- VHDL Architecture DcMotor.valAbsolue.valAbsolue
--
-- Created:
--          by - Aur�lien.UNKNOWN (DESKTOP-24F3HOD)
--          at - 15:53:57 19.08.2019
--
-- using Mentor Graphics HDL Designer(TM) 2015.2 (Build 5)
--
ARCHITECTURE valAbsolue OF valAbsolue IS
BEGIN
END ARCHITECTURE valAbsolue;

