.SUBCKT MCP6547 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following comparators are covered by this model:
*      MCP6546, MCP6547, MCP6548, MCP6549
*
* Revision History:
*      REV A: 16-Oct-07, Created Model
*
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*      Can disable Hysteresis for faster response in large circuits by adding comments
*            in front of statements flagged below
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*      open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit 
*      current, Vsat, Propagation delay vs. Temp and P.S.
*
* Not Supported:
*      Chip Select (MCP6548)
*      Some Variation in specs vs. Power Supply Voltage
*      Monte Carlo (Vos, Ib), Process variation
*      Distortion (detailed non-linear behavior)
*      Behavior outside normal operating region
*
* Input Stage
V10  3 10 -305M
R10 10 11 690K
R11 10 12 690K
G10 10 11 10 11 144U
G11 10 12 10 12 144U
C11 11 12 576E-15
C12  1  0 4P
E12 71 14 POLY(7) 20 0 21 0 22 0 23 0 26 0 27 0 111 0
+ 1.5M 55 55 15 15 1 1 -.5M
* LINE ABOVE FOR HYSTERESIS, LINE BELOW FOR NO HYSTERESIS
*+ 1.5M 55 55 15 15 1 1 0
G12 1 0 62 0 1m
G13 1 2 63 0 1m
M12 11 14 15 15 NMI L=2U W=42U; *Added L & W values
M14 12 2 15 15 NMI L=2U W=42U; *Added L & W values
G14 2 0 62 0 1m
C14  2  0 4P
I15 15 4 50U
I915 4 3 50U
V16 16 4 -305M
GD16 16 1 TABLE {V(16,1)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
V13 3 13 -305M
GD13 2 13 TABLE {V(2,13)} ((-100,-1p)(0,0)(1m,1u)(2m,1m)) 
R71  1  0 20.0E12
R72  2  0 20.0E12
R73  1  2 20.0E12
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G26  0 26 POLY(2) 3 0 4 0   0.00 -160U -160U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -2.75M 133U 133U
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 -2.7
I31 0 31 DC 110
R31 31  0 1 TC=2.34M,-4.57U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 12
I32 32 0 DC 76.5
R32 32  0 1 TC=1.80M,-3.97U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 31.6M
R34  34 0 1K
C34  34 0 503N
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 3P
G38  0 38 37 0 1m
R38  39 0 1K
L38  38 39 32U
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(18.0,1n))(20.0,1))
G36 33 0 TABLE {V(35,4)} ((-22.0,-1)((-20.0,-1n)(0,0)(1,1n))
*
* Output Stage
G57  0 57 POLY(3) 3 0 4 0 35 0   0 -1M -1M -2M
R57 57  4 500
C58  5  0 8P
E58 58 0 VALUE {IF(V(57)>V(3),V(3),IF(V(57)<V(4),V(4),V(57)))}
M5 96 58 4 4 NOUT
*
* Current Limit
R96 96 5 15
D98 4 5 DESD
D99 5 91 DESD
V91 91 4 10
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=2.53M,-13.0U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)} 
+ ((0,0)(600M,5.7N)(650M,30.0N)(800M,200N)
+ (1.33,558N)(1.4,570N)(5.5,580N))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=3.00
E75 1 71 70 0 1 
*
* Temp Sensistive IBias
I62 0 62 DC 1uA
R62 0 62 REXP 68.2U
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1uA
R63 0 63 REXPO 1U
*
* Hysteresis
G110 0 110 POLY(2) 3 0 4 0  3.1 -50M 50M
R110 110 0 1 TC=2.2M,-14U
E111 111 0 VALUE {V(110) * V(112)}
E112 112 0 TABLE {V(120,0)} ((-1,1)(-1m,0.99)(1m,-0.99)(1,-1))
C120  120 0  1u
G120 0 120 TABLE {V(57,4)} ((-1m,-1)(1m,1))
R120 0 120 1
C121 121 120 2p
C122 122 120 2p
V121 121 0 1
V122 122 0 -1
*
* Models
.MODEL NMI NMOS(KP=20U LEVEL=1); *Removed L & W values
.MODEL NOUT NMOS(L=20U W=20U KP=6.7M LEVEL=3 VTO=0.8 VMAX=10000) 
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=146E-18 AF=1
.MODEL REXP  RES TCE= 10.1
.MODEL REXPO RES TCE= 9
.ENDS MCP6547

